module alu (
    input 
);
    
endmodule