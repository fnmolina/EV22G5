module alu (
    input [3:0] operation,
    input [15:0] reg_a, reg_b,
    output reg [3:0] CCR
);
    parameter add = ;
    
endmodule